 -- Illegal Operations 
 JAM_1
 SLO_X_IND
 NOP_ZNG
 SLO_ZPG
 ANC_NUM
 NOP_ABS
 SLO_ABS

 JAM_2
 SLO_IND_Y
 NOP_ZPG_X
 SLO_ZPG_X
 NOP_IMPL
 SLO_ABS_Y
 NOP_ABS_X
 SLO_ABS_X

 JAM_3
 RLA_X_IND
 RLA_ZPG
 ANC_NUM
 RLA_ABS
 
 JAM_4
 RLA_IND_Y
 NOP_ZPG_X
 RLA_ZPG_X
 NOP_IMPL
 RLA_ABS_Y
 NOP_ABS_X
 RLA_ABS_X

 JAM_5
 SRE_X_IND
 NOP_ZPG
 SRE_ZPG
 ALR_NUM
 SRE_ABS

 JAM_6
 SRE_IND_Y
 NOP_ZPG_X
 SRE_ZPG_X
 NOP_IMPL
 SRE_ABS_Y
 NOP_ABS_X
 SRE_ABS_X

 JAM_7
 RRA_X_IND
 NOP_ZPG
 RRA_ZPG
 ARR_NUM
 RRA_ABS

 JAM_8
 RRA_IND_Y
 NOP_ZPG_X
 RRA_ZPG_X
 NOP_IMPL
 RRA_ABS_Y
 NOP_ABS_X
 RRA_ABS_X

 NOP_NUM_1
 NOP_NUM_2
 SAX_X_IND
 SAX_ZPG
 NOP_NUM_3
 ANE_NUM
 SAX_ABS

 JAM_9
 SHA_IND_Y
 SAX_ZPG_Y
 TAS_ABS_Y
 SHA_ABS_X
 SHX_ABS_Y
 SHA_ABS_Y

 LAX_X_IND
 LAX_ZPG
 LXA_NUM
 LAX_ABS

 JAM_10
 LAX_IND_Y
 LAX_ZPG_Y
 LAS_ABS_Y
 LAX_ABS_Y

 NOP_NUM_4
 DCP_X_IND
 DCP_ZPG
 SBX_NUM
 DCP_ABS

 JAM_11
 DCP_IND_Y
 NOP_ZPG_X
 DCP_ZPG_X
 NOP_IMPL
 DCP_ABS_Y
 NOP_ABS_X
 DCP_ABS_X

 NOP_NUM_5
 ISC_X_IND
 ISC_ZPG
 USBC_NUM
 ISC_ABS

 JAM_12
 ISC_IND_Y
 NOP_ZPG_X
 ISC_ZPG_X
 NOP_IMPL
 ISC_ABS_Y
 NOP_ABS_X
 ISC_ABS_X